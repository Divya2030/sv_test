interface mux_if(input logic clk,reset);
  logic sel;
  logic in0;
  logic in1;
  logic out;
endinterface