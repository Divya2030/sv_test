interface count_if(input logic clk,reset);
  logic UpOrDown;
  logic [0:3]count;
endinterface