interface intf_cnt(input logic clk);

    //wire clk;
    logic reset;
    logic data;
    logic [0:3] count;

 endinterface