class scoreboard;
bit  store1;
bit  store2;
bit  store3;
endclass 