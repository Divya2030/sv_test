interface add_if(input logic clk,reset);
  logic a, b,c;
  logic [1:0]sum;
  logic carry;
endinterface