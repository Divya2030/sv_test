 class scoreboard;
       bit  store;
   endclass