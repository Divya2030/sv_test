interface intf_cnt(input logic clk);

    //wire clk;
    logic reset;
    logic din;
    logic dout;

 endinterface